----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/16/2020 04:48:20 PM
-- Design Name: 
-- Module Name: BUFT8 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BUFT8 is
  Port (A : in std_logic_vector (7 downto 0);
        OEn : in std_logic;
        Y : out std_logic_vector (7 downto 0));
end BUFT8;

architecture BUFT8_A of BUFT8 is
begin
    Y <= A when OEn = '0' else "ZZZZZZZZ"; 

end BUFT8_A;
